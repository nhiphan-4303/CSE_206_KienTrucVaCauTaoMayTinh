module Assignment1_Verilog(X,Y,Z);
	input X, Y;
	output Z;
	
	and a1(Z,X,Y);
endmodule